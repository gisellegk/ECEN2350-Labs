/* 
   ECEN 2350: Lab 2
   Module takes number and converts to month and day.  
*/


module dateconverter(input [6:0]num, input leap, output [1:0]month, output [3:0]day_1s, output [1:0]day_10s);
// leap by default is 0 for no leap year. Implement without it for now. 


endmodule